package Basys3Top where

interface Basys3Top =
	-- set leds
	leds :: Bit 16
	-- read switches
	switches :: Bit 16 -> Action
