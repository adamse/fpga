package Basys3Top where

interface SevenSegment =
  seg :: Bit 7
  dp :: Bit 1
  an :: Bit 4

interface Basys3Top =
  buttons :: Buttons
  seven_segment :: SevenSegment
  rs232 :: RS232
  leds :: Bit 16
  switches :: Bit 16 -> Action

interface Buttons =
  bup :: Bool -> Action
  bright :: Bool -> Action
  bdown :: Bool -> Action
  bleft :: Bool -> Action

interface RS232 =
  tx :: Bit 1
  rx :: Bit 1 -> Action
