package Main where

import Vector -- (Vector, (!!), replicate)

import Basys3Top
import ClockDiv

struct ButtonState =
  { up :: Bool
  ; down :: Bool
  ; left :: Bool
  ; right :: Bool
  }
  deriving (Bits)

digitToBits :: UInt 4 -> Bit 7
digitToBits x = case x of
  0 -> 0b1000000
  1 -> 0b1111001
  2 -> 0b0100100
  3 -> 0b0110000
  4 -> 0b0011001
  5 -> 0b0010010
  6 -> 0b0000010
  7 -> 0b1111000
  8 -> 0b0000000
  9 -> 0b0010000
  _ -> 0b1111111

{-# properties mkTop = { alwaysReady, alwaysEnabled } #-}
mkTop :: Module Basys3Top
mkTop = module

  lights_on :: Reg Bool
  lights_on <- mkReg False

  clock :: ClockDiv (UInt 24)
  clock <- mkClockDiv

  switches :: Reg (Bit 16)
  switches <- mkRegU

  pressed_buttons :: Reg ButtonState
  pressed_buttons <- mkReg (ButtonState { up = False; down = False; left = False; right = False })

  seven_segment :: SevenSegment
  seven_segment <- module
    count :: Reg (UInt 4)
    count <- mkReg 0

    pos :: Reg (UInt 2)
    pos <- mkReg 0b00

    rules
      when clock.run_now ==> do
        pos := pos + 1

      when clock.run_now ==> do
        let d =
              if pressed_buttons.up
              then 1
              else if pressed_buttons.down
              then negate 1
              else 0
        count := count + d

    interface
      seg = digitToBits count
      dp = 0b1
      an = case pos of
        0 -> 0b0111
        1 -> 0b1011
        2 -> 0b1101
        3 -> 0b1110

  rules
    when clock.run_now ==> do
      lights_on := not lights_on

  buttons :: Buttons
  buttons <- module
    interface
      bup pressed = pressed_buttons := pressed_buttons { up = pressed }
      bdown pressed = pressed_buttons := pressed_buttons { down = pressed }
      bleft pressed = pressed_buttons := pressed_buttons { left = pressed }
      bright pressed = pressed_buttons := pressed_buttons { right = pressed }

  interface
    leds =
      if lights_on
      then switches
      else 0
    switches values = switches := values
    seven_segment = seven_segment
    buttons = buttons
