module Top (
  output [15:0] led
);

assign led[15] = 1;
assign led[8] = 1;

endmodule
