package Main where

import Clocks

import Basys3Top

struct ButtonState =
  { up :: Reg Bool
  ; down :: Reg Bool
  ; left :: Reg Bool
  ; right :: Reg Bool
  }
  deriving (Bits)

mkButtonState :: Module ButtonState
mkButtonState = module
  up <- mkReg False
  down <- mkReg False
  left <- mkReg False
  right <- mkReg False

  return (ButtonState { up = up; down = down; left = left; right = right })

digitToBits :: UInt 4 -> Bit 7
digitToBits x = case x of
  0 -> 0b1000000
  1 -> 0b1111001
  2 -> 0b0100100
  3 -> 0b0110000
  4 -> 0b0011001
  5 -> 0b0010010
  6 -> 0b0000010
  7 -> 0b1111000
  8 -> 0b0000000
  9 -> 0b0010000
  _ -> 0b1111111

{-# properties mkTop = { alwaysReady, alwaysEnabled } #-}
mkTop :: Module Basys3Top
mkTop = module

  lights_on :: Reg Bool
  lights_on <- mkReg False

  -- 100 mhz default clock
  -- 2 hz
  -- divide by 50m
  two_hz <- mkGatedClockDivider 50_000_000

  switches :: Reg (Bit 16)
  switches <- mkRegU

  pressed_buttons :: ButtonState
  pressed_buttons <- mkButtonState

  seven_segment :: SevenSegment
  seven_segment <- module
    count :: Reg (UInt 4)
    count <- mkReg 0

    pos :: Reg (UInt 2)
    pos <- mkReg 0b00

    rules
      when two_hz.clockReady ==> do
        pos := pos + 1

      when two_hz.clockReady ==> do
        let d =
              if pressed_buttons.up
              then 1
              else if pressed_buttons.down
              then negate 1
              else 0
        count := count + d

    interface
      seg = digitToBits count
      dp = 0b1
      an = case pos of
        0 -> 0b0111
        1 -> 0b1011
        2 -> 0b1101
        3 -> 0b1110

  rules
    when two_hz.clockReady ==> do
      lights_on := not lights_on

  buttons :: Buttons
  buttons <- module
    interface
      bup pressed = pressed_buttons.up := pressed
      bdown pressed = pressed_buttons.down := pressed
      bleft pressed = pressed_buttons.left := pressed
      bright pressed = pressed_buttons.right := pressed

  interface
    leds =
      if lights_on
      then switches
      else 0
    switches values = switches := values
    seven_segment = seven_segment
    buttons = buttons
